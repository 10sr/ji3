module accessmem();
endmodule // accessmem

module alu();